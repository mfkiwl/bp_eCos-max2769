# ====================================================================
#
#      ser_arm_bp2016.cdl
#
#      eCos serial ARM/BP2016 configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      michael anburaj <michaelanburaj@hotmail.com>
# Contributors:   michael anburaj <michaelanburaj@hotmail.com>
# Date:           2003-08-01
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_ARM_BP2016 {
    display       "HG BP2016 board serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_ARM_BP2016

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    include_files ; # none _exported_ whatsoever
    description   "
           This option enables the serial device drivers for the
           HG BP2016 based development boards."

    compile       -library=libextras.a   bp2016_serial.c uart_api.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_arm_bp2016.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_BP2016_UART_FIFO {
        display       "bp2016 FIFO support"
        flavor        bool
        default_value 1
        description   "
            Options to configure the FIFO on bp2016."
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL0 {
        display       "HG BP2016 serial port 0 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for the HG BP2016 port 0."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL0_NAME {
            display       "Device name for the HG BP2016 serial port 0 driver"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL0_BAUD {
            display       "Baud rate for the HG BP2016 serial port 0 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL0_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 0 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 256
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL0_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 0 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 0."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL0_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL0_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL0_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 0 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 0."
        }
	}

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL1 {
        display       "HG BP2016 serial port 1 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the HG BP2016 port 1."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL1_NAME {
            display       "Device name for the HG BP2016 serial port 1 driver"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL1_BAUD {
            display       "Baud rate for the HG BP2016 serial port 1 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL1_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 1 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 8192
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL1_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 1 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 1."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL1_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL1_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL1_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 1 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 1."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL2 {
        display       "HG BP2016 serial port 2 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the HG BP2016 port 2."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL2_NAME {
            display       "Device name for the HG BP2016 serial port 2 driver"
            flavor        data
            default_value {"\"/dev/ser2\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 2."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL2_BAUD {
            display       "Baud rate for the HG BP2016 serial port 2 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 2."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL2_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 2 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 256
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 2."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL2_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 2 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 2."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL2_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL2_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL2_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 1 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 2."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL3 {
        display       "HG BP2016 serial port 3 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the HG BP2016 port 3."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL3_NAME {
            display       "Device name for the HG BP2016 serial port 3 driver"
            flavor        data
            default_value {"\"/dev/ser3\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 3."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL3_BAUD {
            display       "Baud rate for the HG BP2016 serial port 3 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 3."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL3_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 3 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 256
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 3."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL3_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 3 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 3."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL3_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL3_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL3_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 3 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 3."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL4 {
        display       "HG BP2016 serial port 4 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the HG BP2016 port 4."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL4_NAME {
            display       "Device name for the HG BP2016 serial port 4 driver"
            flavor        data
            default_value {"\"/dev/ser4\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 4."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL4_BAUD {
            display       "Baud rate for the HG BP2016 serial port 4 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 4."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL4_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 4 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 256
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 4."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL4_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 4 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 4."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL4_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL4_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL4_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 4 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 4."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL5 {
        display       "HG BP2016 serial port 5 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for the HG BP2016 port 5."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL5_NAME {
            display       "Device name for the HG BP2016 serial port 5 driver"
            flavor        data
            default_value {"\"/dev/ser5\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 5."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL5_BAUD {
            display       "Baud rate for the HG BP2016 serial port 5 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 5."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL5_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 5 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 256
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 5."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL5_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 1 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 5."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL5_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL5_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL5_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 1 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 5."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL6 {
        display       "HG BP2016 serial port 6 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for the HG BP2016 port 6."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL6_NAME {
            display       "Device name for the HG BP2016 serial port 6 driver"
            flavor        data
            default_value {"\"/dev/ser6\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 6."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL6_BAUD {
            display       "Baud rate for the HG BP2016 serial port 6 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
                          460800 921600 1875000 2850000
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 6."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL6_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 6 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 8192
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 6."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL6_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 6 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 6."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL6_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL6_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL6_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 6 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 6."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_SERIAL7 {
        display       "HG BP2016 serial port 7 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for the HG BP2016 port 7."

        cdl_option CYGDAT_IO_SERIAL_ARM_BP2016_SERIAL7_NAME {
            display       "Device name for the HG BP2016 serial port 7 driver"
            flavor        data
            default_value {"\"/dev/ser7\""}
            description   "
                This option specifies the name of serial device for the HG BP2016 port 7."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL7_BAUD {
            display       "Baud rate for the HG BP2016 serial port 7 driver"
            flavor        data
            legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                          4800 7200 9600 14400 19200 38400 57600 115200 230400
                          460800 921600 1875000 2850000
            }
            default_value 115200
            description   "
                This option specifies the default baud rate (speed) for the HG BP2016 port 7."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL7_BUFSIZE {
            display       "Buffer size for the HG BP2016 serial port 7 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 8192
            description   "
                This option specifies the size of the internal buffers used for
                the HG BP2016 port 7."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL7_FIFOSIZE {
            display       "Buffer size for the HG BP2016 serial port 7 driver"
            flavor        data
            legal_values  256
            default_value 256
            description   "
                This option specifies the size of the hardware fifo used for
                the HG BP2016 port 7."
        }

        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL7_FIFO_RX_THRESHOLD {
            display "Threshold for RX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the RX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--1 character in fifo,
                1--1/4 full of fifo,
                2--1/2 of fifo depth,
                3--2 less than full."
        }
        cdl_option CYGPKG_IO_SERIAL_BP2016_SERIAL7_FIFO_TX_THRESHOLD {
            display "Threshold for TX interrupt on 16550 FIFO"
            flavor data
            legal_values { 3 2 1 0 }
            default_value 0
            description "
                This options configures the threshold value at which
                the TX interrupt occurs when a FIFO is used. (16550 and
                above only)
                0--acturally empty,
                1--2 characters left in tx fifo,
                2--1/4 of fifo depth,
                3--1/2 of fifo depth."
        }

        cdl_option CYGNUM_IO_SERIAL_ARM_BP2016_SERIAL7_AUTO_FLOW_CONTROL {
            display       "Auto flow control for the HG BP2016 serial port 1 driver"
            flavor data
            legal_values { 1 0 }
            default_value 0
            description   "
                This option specifies the auto flow control enable status for
                the HG BP2016 port 7."
        }
    }


    cdl_component CYGPKG_IO_SERIAL_ARM_BP2016_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
            Package specific build options including control over
            compiler flags used only in building this package,
            and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_ARM_BP2016_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_ARM_BP2016_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

}

# EOF ser_arm_bp2016.cdl
