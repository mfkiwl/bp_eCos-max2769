# ====================================================================
#
#      hal_arm_bp2016_asic.cdl
#
#      HG BP2016 asic package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2006 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Mike Jones
# Contributors:
# Date:           2013-08-08
#
#####DESCRIPTIONEND####

cdl_package CYGPKG_HAL_ARM_BP2016_ASIC_BP_SIDE {

    display       "HG BP2016 ASIC board"
    parent         CYGPKG_HAL_ARM_BP2016

    include_dir    cyg/hal
    define_header  hal_arm_bp2016_asic.h
    hardware

    description    "
        This HAL platform package provides generic
        support for the bp2016 asic board."

    compile       asic_misc.c platform_init.c 

    implements    CYGINT_HAL_ARM_ARCH_ARM_CORTEXA7

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_bp2016.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_bp2016_asic.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"Cortex-A7\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"BP2016 ASIC\""
    }

    cdl_option CYGHWR_HAL_BP2016_SUPPORT_FAST_BOOT {
        display          "Enable Fast booting for BP side"
        default_value    0
        description      "
            Enable Fast booting."
    }

    cdl_option CYGHAL_RUN_ENV_DDR {
        display       "Running on ddr or not"
            flavor        bool
            default_value 0
            description   "Select firmware running on ddr or not"
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { (CYG_HAL_STARTUP == "RAM") ? "arm_asic_ram" : "arm_asic_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { (CYGHAL_RUN_ENV_DDR == 1) ? "<pkgconf/mlt_arm_asic_ddr.ldi>" : "<pkgconf/mlt_arm_asic_ram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { (CYGHAL_RUN_ENV_DDR == 1) ? "<pkgconf/mlt_arm_asic_ddr.h>" : "<pkgconf/mlt_arm_asic_ram.h>" }
        }
    }
    cdl_option CYGNUM_HAL_RTC_TIMER_ID {
        display          "RTC Timer id"
        flavor data
        legal_values     0 to 3
        default_value    0
        description      "
            The asic has 4 ext-timer. This option
            chooses which timer will be used to os tick."
     }
    
    cdl_option CYGNUM_HAL_KERNEL_COUNTERS_CLOCK_ISR_DEFAULT_PRIORITY {
	    display		"Default priority for system clock interrupts"
	    flavor		data
        default_value 160
	    description "
            The Bp2016 eCos HAL RTC priority Default value."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display       "Number of communication channels on the board"
        flavor        data
        calculated    8
        description   "
            The Evk board has one serial port: UART0."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The asic has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The asic board has two UART serial ports. This option
            chooses which port will be used for diagnostic output."
     }
     
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the diagnostic port."
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
         display       "GDB serial port baud rate"
         flavor        data
         legal_values  9600 19200 38400 57600 115200
         default_value 115200 
         description   "
            This option controls the baud rate used for the GDB connection."
     }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . CYGBLD_ARCH_CFLAGS .
                            "-Wstrict-prototypes -Wno-comment -mcpu=cortex-a7 -mfloat-abi=softfp -mfpu=neon -g -Os -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -ffreestanding" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGBLD_ARCH_LDFLAGS . "-mcpu=cortex-a7 -static -n -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

}
#-mfloat-abi=hard 
