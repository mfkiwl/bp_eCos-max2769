# ====================================================================
#
#      hal_arm_bp2016.cdl
#
#      HG BP2016 HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      zhijiehao
# Contributors:   
# Date:           2017-01-18
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_BP2016 {
    display       "HG BP2016 variant HAL"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_bp2016.h
    include_dir   cyg/hal
    hardware
    description   "
        The bp2016 HAL package provides the support needed to run
        eCos on HG bp2016 based targets."

    compile		bp2016_timer.c bp2016_intr.c bp2016_plf_misc.c bp2016_scm.c bp2016_gpio.c timer/timer_imp.c uart/uart_imp.c gic/gic400.c a7/cache_v7.c a7/mmu_setup.c a7/arch_timer.c a7/v7_cp15.S a7/memcpy.S a7/memset.S sim/sim.c sim/sim_hal.c clk/clk_hw.c reset/reset_hw.c  gpio/gpio_imp.c spi/spi_dw.c spi/spi3wire.c gpio/gpio_api.c dma/dma_imp.c backtrace/backtrace.c misc/wakeupap.c
	compile		iomux/iomux_hw_gpio.c iomux/iomux_hw_mmc.c iomux/iomux_hw_pwm.c iomux/iomux_hw_sim.c iomux/iomux_hw_sram.c iomux/iomux_hw_if.c iomux/iomux_hw_prm.c iomux/iomux_hw_regs.c iomux/iomux_hw_scm.c iomux/iomux_hw_spi.c iomux/iomux_hw_uart.c iomux/iomux_hw_api.c
	compile		backtrace/dump_stack.c misc/debug_misc.c
	compile		comm/cpu_comm.c
	compile		asram/asram.c
	compile		misc/rsv_data.c
    compile     wdt/wdt_hw.c wdt/wdt_api.c 
    compile     pll/pll.c pll/pll_api.c 
    compile     gpio/spi4_bitbang.c
    compile     gpio/spi_bitbang.c
    compile     pwm/pwm.c pwm/pwm_api.c
    compile     misc/fastboot_reset.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT
    implements    CYGINT_HAL_ARM_ARCH_ARM_CORTEXA7
    implements    CYGINT_HAL_ARM_THUMB_ARCH
    #requires      CYGDBG_USE_ASSERTS
    #requires      CYGIMP_KERNEL_SCHED_SORTED_QUEUES

	cdl_option CYGFUN_KERNEL_THREADS_SWITCH_STATS {
        display    "thread switches statistics support"
        calculated 0
        description    "thread switches statistics support."
    }

	cdl_component CYGNUM_KERNEL_TREAHD_STATS {
        display        "statistics thread max number"
        flavor         data
        default_value  32
        description "statistics thread max number"
    }

    cdl_option CYGHWR_HAL_ARM_FPU {
        display    "Variant FPU support"
        calculated 1
        description    "The bp2016 supports VFPv4 instructions."
    }

    cdl_option CYGHWR_HAL_ARM_FPU_D32 {
        display    "Variant vfpvxu-d32 support"
        calculated 1
        description    "The bp2016 supports VFPv4-d32 instructions."
    }


    cdl_option CYGHWR_HAL_ARM_NEON {
        display    "Variant NEON support"
        calculated 1
        description    "The bp2016 supports NEON instructions."
    }

    # Let the architectural HAL see this variant's files
    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_ARCH_H"
    }

    cdl_option CYGHWR_HAL_ARM_BP2016 {
        display        "BP2016 variant used"
        flavor         data
        default_value  {"BP2016UL"}
        legal_values   {"BP2016UL"}
        description    "The bp2016 microcontroller family has several variants,
			This option allows the platform HALs to select the 
                        specific microcontroller being used."
    }

    cdl_option CYGINT_HAL_INTERRUPT_TIME_STAT {
	    display     "Platform provides the time statistics for per irq"
        calculated 1
	    description "Only for debug function, when debug system performance"
    }


    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "Norflash" }
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            When targeting the bp2016 eval boards it is only possible to build
            the system for RAM bootstrap."
    }

    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
               
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
	    calculated    950000
            description   "Value to program into the RTC clock generator. OS timer must be 10 ms."
        }
    }

    cdl_component CYGNUM_HAL_STARTUP_STACK_SIZE {
        display        "Starutp stack size"
        flavor         data
        default_value  2048
        description "
            Size of the startup stack used during initialization
             of the system."
    }

    cdl_component CYGDBG_RELEASE_MSG {
        display        "Release message"
        flavor         data
        default_value  1
        description "release message."

    cdl_option CYGDBG_RELEASE_VERSION {
        display        "release version"
        flavor         data
        default_value  170
        description "release version."
    }

    cdl_option CYGDBG_RELEASE_TYPE {
        display        "release type"
        flavor         data
        default_value  { 0 }
        legal_values   { 0 1 }
        description    "
                        this is choise for cpu0 or cpu1."
    }

    cdl_option CYGHWR_HAL_ASIC_CLK {
        display        "bp2016 asic contains clock settings"
        flavor         bool
        default_value  { 0 }
    }

	make -priority 50 {
	    <PREFIX>/include/cyg/hal/version.h: <PACKAGE>/cdl/hal_arm_bp2016.cdl
	    sh $(REPOSITORY)/$(PACKAGE)/script/version.sh $< > $@
	}
    }
}
